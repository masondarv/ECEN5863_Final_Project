// Doty Darveaux
// ECEN 5863
// Pong Final Project

module collision(
	input clk, reset,
	input paddle_1_sig,
	input paddle_2_sig,
	input ball_sig,
	input frame_sig,
	output collision);

endmodule // frame