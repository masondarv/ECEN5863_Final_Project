
module paddle(
input clk, rst,
input [9:0] hcount, vcount,
output r, g, b
);


endmodule
