// Doty Darveaux
// ECEN 5863
// Pong Final Project

module collision(
	input clk, reset,
	input paddle_1_r, paddle_1_g, paddle_1_b,
	input paddle_2_r, paddle_2_g, paddle_2_b,
	input ball_r, ball_g, ball_b,
	input frame_r, frame_g, frame_b,
	output r, g, b );

endmodule // frame