// Doty Darveaux
// ECEN 5863
// Pong Final Project

module frame(
	input clk, reset,
	input [9:0] hcount, vcount,
	output r, g, b );

endmodule // frame